// 2016 Ryan Leonard
// RegisterFile (RF) Module Testbench

module rf_32_test
