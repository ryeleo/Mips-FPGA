// 2016 Ryan Leonard
// RegisterFile (RF) Module Testbench

module registerFile_test
